magic
tech sky130A
magscale 1 2
timestamp 1680637778
<< nwell >>
rect 7076 -1112 7446 250
<< locali >>
rect 194 940 8090 976
rect 194 842 506 940
rect 8028 842 8090 940
rect 194 820 8090 842
rect 190 726 8090 820
rect 190 -408 1182 726
rect 190 -956 350 -408
rect 814 -956 1182 -408
rect 184 -1606 366 -1172
rect 1704 -1182 2076 726
rect 2810 -1176 3182 726
rect 4540 222 8090 726
rect 4540 164 8088 222
rect 4540 18 7446 164
rect 4540 -1168 4912 18
rect 7076 -1112 7446 18
rect 7764 -1102 8088 164
rect 848 -1432 8080 -1316
rect 834 -1476 8080 -1432
rect 184 -1610 654 -1606
rect 834 -1610 2766 -1476
rect 184 -1712 2766 -1610
rect 184 -1796 2608 -1712
rect 184 -2176 654 -1796
rect 2552 -2176 2608 -1796
rect 184 -2238 2608 -2176
rect 2730 -2176 2766 -1712
rect 7116 -1710 8074 -1476
rect 7116 -2176 7198 -1710
rect 2730 -2234 7198 -2176
rect 7302 -1842 8074 -1710
rect 7302 -2176 7424 -1842
rect 7750 -2176 8074 -1842
rect 7302 -2234 8080 -2176
rect 2730 -2238 8080 -2234
rect 184 -2288 8080 -2238
rect 184 -2386 440 -2288
rect 7974 -2386 8080 -2288
rect 184 -2426 8080 -2386
<< viali >>
rect 506 842 8028 940
rect 2608 -2238 2730 -1712
rect 7198 -2234 7302 -1710
rect 440 -2386 7974 -2288
<< metal1 >>
rect 186 940 8080 978
rect 186 842 506 940
rect 8028 842 8080 940
rect 186 740 8080 842
rect 1358 608 1562 740
rect 1226 134 1236 458
rect 1302 134 1312 458
rect 1588 134 1598 458
rect 1664 134 1674 458
rect 194 -286 620 -40
rect 384 -1064 448 -602
rect 368 -1194 378 -1064
rect 450 -1194 460 -1064
rect 384 -1448 448 -1194
rect 550 -1518 616 -286
rect 693 -743 1008 -657
rect 922 -1038 1008 -743
rect 922 -1124 1542 -1038
rect 724 -2032 776 -1364
rect 1826 -2104 1966 740
rect 2244 624 2644 740
rect 3322 634 3332 690
rect 3704 634 3714 690
rect 4008 634 4018 690
rect 4390 634 4400 690
rect 2114 136 2124 456
rect 2200 136 2210 456
rect 2682 132 2692 452
rect 2768 132 2778 452
rect 2246 -632 2644 -616
rect 2246 -920 2262 -632
rect 2626 -920 2644 -632
rect 2246 -1060 2644 -920
rect 3240 -930 3250 -620
rect 3304 -930 3314 -620
rect 3432 -1066 3594 634
rect 3752 -1070 3846 602
rect 3926 -930 3936 -620
rect 3990 -930 4000 -620
rect 4116 -1060 4278 634
rect 3740 -1196 3750 -1070
rect 3852 -1196 3862 -1070
rect 3752 -1504 3846 -1196
rect 4444 -1324 4552 602
rect 7566 434 7644 448
rect 7204 422 7256 428
rect 7204 364 7256 370
rect 5058 2 6928 4
rect 4962 -66 6928 2
rect 4962 -90 5088 -66
rect 4962 -208 5088 -194
rect 4960 -440 4970 -208
rect 5040 -440 5088 -208
rect 4962 -446 5088 -440
rect 5292 -1000 5570 -66
rect 5842 -70 5950 -66
rect 5840 -92 5950 -70
rect 5862 -162 5950 -92
rect 5374 -1066 5542 -1060
rect 5362 -1200 5372 -1066
rect 5542 -1200 5552 -1066
rect 4432 -1432 4442 -1324
rect 4550 -1432 4560 -1324
rect 4840 -1328 4948 -1318
rect 4828 -1436 4838 -1328
rect 4946 -1436 4956 -1328
rect 4840 -1504 4948 -1436
rect 2918 -1600 3846 -1504
rect 4000 -1600 4948 -1504
rect 2592 -1696 2750 -1688
rect 2434 -2186 2512 -1952
rect 2588 -1968 2598 -1696
rect 2746 -1968 2756 -1696
rect 2830 -1968 2840 -1700
rect 2902 -1968 2912 -1700
rect 2592 -2186 2608 -1968
rect 186 -2238 2608 -2186
rect 2730 -2186 2750 -1968
rect 3230 -2096 3396 -1600
rect 3752 -2032 3846 -1600
rect 3916 -1970 3926 -1702
rect 3988 -1970 3998 -1702
rect 4328 -2098 4494 -1600
rect 4840 -2056 4948 -1600
rect 5004 -1968 5014 -1700
rect 5076 -1968 5086 -1700
rect 5374 -2098 5542 -1200
rect 5896 -1222 5950 -162
rect 6046 -444 6056 -212
rect 6126 -444 6136 -212
rect 6400 -998 6678 -66
rect 6988 -144 7102 -130
rect 6970 -1176 7102 -144
rect 5896 -1276 5991 -1222
rect 5937 -2045 5991 -1276
rect 6480 -1432 6490 -1326
rect 6640 -1432 6650 -1326
rect 6090 -1970 6100 -1702
rect 6162 -1970 6172 -1702
rect 6480 -2098 6648 -1432
rect 6962 -1500 6972 -1176
rect 7048 -1490 7102 -1176
rect 7208 -1478 7252 364
rect 7556 180 7566 434
rect 7648 180 7658 434
rect 7574 42 7640 180
rect 7794 -8 7998 740
rect 7510 -444 7520 -210
rect 7578 -444 7588 -210
rect 7646 -986 7998 -8
rect 7646 -1218 7762 -1206
rect 7646 -1478 7660 -1218
rect 7748 -1478 7762 -1218
rect 7048 -1500 7082 -1490
rect 6992 -1510 7082 -1500
rect 6998 -1648 7082 -1510
rect 7208 -1518 7604 -1478
rect 7208 -1520 7252 -1518
rect 6992 -2038 7082 -1648
rect 7180 -1698 7312 -1696
rect 7170 -1968 7180 -1698
rect 7314 -1968 7324 -1698
rect 6514 -2108 6622 -2098
rect 7180 -2186 7198 -1968
rect 2730 -2234 7198 -2186
rect 7302 -2186 7312 -1968
rect 7564 -1976 7604 -1518
rect 7478 -2186 7558 -2008
rect 7646 -2106 7762 -1478
rect 7302 -2234 8080 -2186
rect 2730 -2238 8080 -2234
rect 186 -2288 8080 -2238
rect 186 -2386 440 -2288
rect 7974 -2386 8080 -2288
rect 186 -2424 8080 -2386
<< via1 >>
rect 1236 134 1302 458
rect 1598 134 1664 458
rect 378 -1194 450 -1064
rect 3332 634 3704 690
rect 4018 634 4390 690
rect 2124 136 2200 456
rect 2692 132 2768 452
rect 2262 -920 2626 -632
rect 3250 -930 3304 -620
rect 3936 -930 3990 -620
rect 3750 -1196 3852 -1070
rect 7204 370 7256 422
rect 4970 -440 5040 -208
rect 5372 -1200 5542 -1066
rect 4442 -1432 4550 -1324
rect 4838 -1436 4946 -1328
rect 2598 -1712 2746 -1696
rect 2598 -1968 2608 -1712
rect 2608 -1968 2730 -1712
rect 2730 -1968 2746 -1712
rect 2840 -1968 2902 -1700
rect 3926 -1970 3988 -1702
rect 5014 -1968 5076 -1700
rect 6056 -444 6126 -212
rect 6490 -1432 6640 -1326
rect 6100 -1970 6162 -1702
rect 6972 -1500 7048 -1176
rect 7566 180 7648 434
rect 7520 -444 7578 -210
rect 7660 -1478 7748 -1218
rect 7180 -1710 7314 -1698
rect 7180 -1968 7198 -1710
rect 7198 -1968 7302 -1710
rect 7302 -1968 7314 -1710
<< metal2 >>
rect 3398 700 3664 1228
rect 4068 700 4334 1228
rect 3332 690 3704 700
rect 3332 624 3704 634
rect 4018 690 4390 700
rect 4018 624 4390 634
rect 1236 458 1302 468
rect 1598 458 1664 468
rect 2124 458 2200 466
rect 2692 458 2768 462
rect 182 134 1236 458
rect 1302 134 1598 458
rect 1664 456 2768 458
rect 1664 136 2124 456
rect 2200 452 2768 456
rect 2200 136 2692 452
rect 1664 134 2692 136
rect 1236 124 1302 134
rect 1598 124 1664 134
rect 2124 126 2200 134
rect 7566 434 7648 444
rect 2768 422 7566 430
rect 2768 370 7204 422
rect 7256 370 7566 422
rect 2768 180 7566 370
rect 7648 180 7654 430
rect 2768 178 7654 180
rect 7566 170 7648 178
rect 2692 122 2768 132
rect 4970 -208 5040 -198
rect 6056 -208 6126 -202
rect 7520 -208 7578 -200
rect 5040 -210 7590 -208
rect 5040 -212 7520 -210
rect 5040 -440 6056 -212
rect 4970 -442 6056 -440
rect 4970 -450 5040 -442
rect 6126 -442 7520 -212
rect 6056 -454 6126 -444
rect 7578 -442 7590 -210
rect 7520 -454 7578 -444
rect 3250 -616 3304 -610
rect 3936 -616 3990 -610
rect 2128 -620 4522 -616
rect 2128 -632 3250 -620
rect 2128 -920 2262 -632
rect 2626 -920 3250 -632
rect 2128 -930 3250 -920
rect 3304 -930 3936 -620
rect 3990 -930 4522 -620
rect 2128 -934 4522 -930
rect 3250 -940 3304 -934
rect 3936 -940 3990 -934
rect 378 -1064 450 -1054
rect 3750 -1068 3852 -1060
rect 5372 -1066 5542 -1056
rect 450 -1070 5372 -1068
rect 450 -1194 3750 -1070
rect 378 -1196 3750 -1194
rect 3852 -1196 5372 -1070
rect 378 -1204 450 -1196
rect 3750 -1206 3852 -1196
rect 5542 -1196 5644 -1068
rect 6972 -1174 7048 -1166
rect 6972 -1176 8072 -1174
rect 5372 -1210 5542 -1200
rect 4442 -1324 4550 -1314
rect 4838 -1324 4946 -1318
rect 6490 -1324 6640 -1316
rect 4550 -1326 6640 -1324
rect 4550 -1328 6490 -1326
rect 4550 -1432 4838 -1328
rect 4442 -1442 4550 -1432
rect 4946 -1432 6490 -1328
rect 4838 -1446 4946 -1436
rect 6490 -1442 6640 -1432
rect 7048 -1218 8072 -1176
rect 7048 -1478 7660 -1218
rect 7748 -1478 8072 -1218
rect 7048 -1500 8072 -1478
rect 6972 -1510 7048 -1500
rect 2598 -1696 2746 -1686
rect 2840 -1696 2902 -1690
rect 3926 -1696 3988 -1692
rect 5014 -1696 5076 -1690
rect 6100 -1696 6162 -1692
rect 7180 -1696 7314 -1688
rect 2746 -1698 7314 -1696
rect 2746 -1700 7180 -1698
rect 2746 -1968 2840 -1700
rect 2902 -1702 5014 -1700
rect 2902 -1968 3926 -1702
rect 2598 -1970 3926 -1968
rect 3988 -1968 5014 -1702
rect 5076 -1702 7180 -1700
rect 5076 -1968 6100 -1702
rect 3988 -1970 6100 -1968
rect 6162 -1968 7180 -1702
rect 6162 -1970 7314 -1968
rect 2598 -1978 2746 -1970
rect 2840 -1978 2902 -1970
rect 3926 -1980 3988 -1970
rect 5014 -1978 5076 -1970
rect 6100 -1980 6162 -1970
rect 7180 -1978 7314 -1970
use sky130_fd_pr__pfet_01v8_GGMWVD  XM1
timestamp 1680634426
transform 0 1 1449 -1 0 -200
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM2
timestamp 1680634426
transform 1 0 3316 0 1 -1840
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM3
timestamp 1680634426
transform 1 0 3516 0 1 -195
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_GGY9VD  XM4
timestamp 1680634426
transform 0 1 2441 -1 0 -204
box -996 -419 996 419
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM5
timestamp 1680634426
transform 1 0 6542 0 1 -531
box -596 -619 596 619
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM6
timestamp 1680634426
transform 1 0 6574 0 1 -1840
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_L9KS9E  XM7
timestamp 1680636816
transform 1 0 7585 0 1 -2031
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM8
timestamp 1680634426
transform 1 0 574 0 1 -677
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_lvt_FMMQLY  XM9
timestamp 1680634426
transform 1 0 598 0 1 -1402
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_lvt_FMHZDY  XM10
timestamp 1680634426
transform 1 0 1606 0 1 -1996
box -996 -260 996 260
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM12
timestamp 1680634426
transform 1 0 5488 0 1 -1840
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM18
timestamp 1680634426
transform 1 0 4402 0 1 -1840
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM20
timestamp 1680634426
transform 1 0 4202 0 1 -195
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_MGSVTJ  XM46
timestamp 1680636816
transform 1 0 7607 0 1 -464
box -211 -684 211 684
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM54
timestamp 1680634426
transform 1 0 5456 0 1 -531
box -596 -619 596 619
<< labels >>
flabel metal1 220 762 420 962 0 FreeSans 256 0 0 0 VCC
port 5 nsew
flabel metal1 216 -2394 416 -2194 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal2 3426 1002 3626 1202 0 FreeSans 256 0 0 0 MINUS
port 2 nsew default input
flabel metal2 4112 1002 4312 1202 0 FreeSans 256 0 0 0 PLUS
port 1 nsew default input
flabel metal2 230 212 430 412 0 FreeSans 256 0 0 0 EN_N
port 3 nsew
flabel metal2 7840 -1430 8040 -1230 0 FreeSans 256 0 0 0 DIFFOUT
port 6 nsew
flabel metal1 214 -266 414 -66 0 FreeSans 256 0 0 0 ADJ
port 7 nsew
flabel metal2 2982 -792 2982 -792 0 FreeSans 800 0 0 0 SP
flabel metal1 3796 -1298 3796 -1298 0 FreeSans 800 0 0 0 G1
flabel metal1 4498 -1250 4498 -1250 0 FreeSans 800 0 0 0 G2
<< end >>
