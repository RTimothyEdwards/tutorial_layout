magic
tech sky130A
magscale 1 2
timestamp 1680636816
<< error_p >>
rect -29 545 29 551
rect -29 511 -17 545
rect -29 505 29 511
<< nwell >>
rect -211 -684 211 684
<< pmos >>
rect -15 -536 15 464
<< pdiff >>
rect -73 452 -15 464
rect -73 -524 -61 452
rect -27 -524 -15 452
rect -73 -536 -15 -524
rect 15 452 73 464
rect 15 -524 27 452
rect 61 -524 73 452
rect 15 -536 73 -524
<< pdiffc >>
rect -61 -524 -27 452
rect 27 -524 61 452
<< nsubdiff >>
rect -175 614 -79 648
rect 79 614 175 648
rect -175 551 -141 614
rect 141 551 175 614
rect -175 -614 -141 -551
rect 141 -614 175 -551
rect -175 -648 -79 -614
rect 79 -648 175 -614
<< nsubdiffcont >>
rect -79 614 79 648
rect -175 -551 -141 551
rect 141 -551 175 551
rect -79 -648 79 -614
<< poly >>
rect -33 545 33 561
rect -33 511 -17 545
rect 17 511 33 545
rect -33 495 33 511
rect -15 464 15 495
rect -15 -562 15 -536
<< polycont >>
rect -17 511 17 545
<< locali >>
rect -175 614 -79 648
rect 79 614 175 648
rect -175 551 -141 614
rect 141 551 175 614
rect -33 511 -17 545
rect 17 511 33 545
rect -61 452 -27 468
rect -61 -540 -27 -524
rect 27 452 61 468
rect 27 -540 61 -524
rect -175 -614 -141 -551
rect 141 -614 175 -551
rect -175 -648 -79 -614
rect 79 -648 175 -614
<< viali >>
rect -17 511 17 545
rect -61 -524 -27 452
rect 27 -524 61 452
<< metal1 >>
rect -29 545 29 551
rect -29 511 -17 545
rect 17 511 29 545
rect -29 505 29 511
rect -67 452 -21 464
rect -67 -524 -61 452
rect -27 -524 -21 452
rect -67 -536 -21 -524
rect 21 452 67 464
rect 21 -524 27 452
rect 61 -524 67 452
rect 21 -536 67 -524
<< properties >>
string FIXED_BBOX -158 -631 158 631
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
